module m310_hpec_subsys_main(
	input aaa;
	input bbb;
	
	output ccc;
	output [31:0] ddd;

);
assign ccc = 0;
assign ddd[31:0]  = 0;
endmodule
